typedef uvm_reg_field rggen_ral_field;
