class rggen_ral_field extends rggen_ral_field_base;
  function new(string name = "rggen_ral_field");
    super.new(name);
  endfunction
endclass
