class rggen_ral_block extends uvm_reg_block;
  function new(string name, int has_coverage = UVM_NO_COVERAGE);
    super.new(name, has_coverage);
  endfunction

  function void configure(
    uvm_reg_block parent    = null,
    string        hdl_path  = ""
  );
    super.configure(parent, hdl_path);
    if (default_map == null) begin
      default_map = create_default_map();
    end
  endfunction

  function void lock_model();
    uvm_reg_block parent;
    uvm_reg_map   maps[$];

    if (is_locked()) begin
      return;
    end

    super.lock_model();
    parent  = get_parent();
    if (parent != null) begin
      return;
    end

    get_maps(maps);
    foreach (maps[i]) begin
      rggen_ral_map rggen_map;
      if ($cast(rggen_map, maps[i])) begin
        rggen_map.Xinit_indirect_reg_address_mapX();
      end
    end
  endfunction

  virtual function uvm_reg_map create_map(
    string            name,
    uvm_reg_addr_t    base_addr,
    int unsigned      n_bytes,
    uvm_endianness_e  endian,
    bit               byte_addressing = 1
  );
    uvm_factory f = uvm_factory::get();
    f.set_inst_override_by_type(
      uvm_reg_map::get_type(), rggen_ral_map::get_type(), {get_full_name(), ".", name}
    );
    return super.create_map(name, base_addr, n_bytes, endian, byte_addressing);
  endfunction

  protected virtual function uvm_reg_map create_default_map();
    return null;
  endfunction
endclass
