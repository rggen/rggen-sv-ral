class rggen_ral_reg_file extends rggen_ral_block;
  protected int unsigned  array_index[$];

  function new(string name, int unsigned n_bytes);
    super.new(name, n_bytes);
  endfunction

  function void configure(
    uvm_reg_block parent,
    int unsigned  array_index[$],
    string        hdl_path
  );
    super.configure(parent, hdl_path);
    foreach (array_index[i]) begin
      this.array_index.push_back(array_index[i]);
    end
  endfunction

  virtual function rggen_ral_block get_block();
    rggen_ral_reg_file  file;
    rggen_ral_block     block;

    if ($cast(file, get_parent())) begin
      return file.get_parent();
    end
    else if ($cast(block, get_parent())) begin
      return block;
    end
    else begin
      return null;
    end
  endfunction

  virtual function void get_array_index(ref int unsigned array_index[$]);
    foreach (this.array_index[i]) begin
      array_index.push_back(this.array_index[i]);
    end
  endfunction
endclass
